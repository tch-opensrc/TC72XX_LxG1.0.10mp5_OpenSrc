PO4A-HEADER:mode=after;position=F�RFATTARE;beginboundary=.SH
.SH �VERS�TTNING
David Weinehall
.RI < tao@kernel.org >
